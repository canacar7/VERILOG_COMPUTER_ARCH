`timescale 1ns / 1ps

module mux4x32_tb();
	
	reg [31 : 0] a0,a1,a2,a3;
	reg  [1: 0]  s;
	wire [31: 0] y;
	
	mux4x32 m_aktif(a0,a1,a2,a3,s,y);
	
	initial begin
	
		#5 a0 = 32'hF0000000; a1 = 32'h00000000; a2 = 32'hF0000000; a3 = 32'h00000000;  s = 00;
		#5 a0 = 32'hF0000001; a1 = 32'h00000001; a2 = 32'hF0000001; a3 = 32'h00000001;  s = 01;
		#5 a0 = 32'hF0000010; a1 = 32'h00000010; a2 = 32'hF0000010; a3 = 32'h00000010;  s = 00;
		#5 a0 = 32'hF0000100; a1 = 32'h00000100; a2 = 32'hF0000100; a3 = 32'h00000100;  s = 01;
		#5 a0 = 32'hF0001000; a1 = 32'h00001000; a2 = 32'hF0001000; a3 = 32'h00001000;  s = 00;
		#5 a0 = 32'hF0010000; a1 = 32'h00010000; a2 = 32'hF0010000; a3 = 32'h00010000;  s = 00;
		#5 a0 = 32'hF0100000; a1 = 32'h00100000; a2 = 32'hF0100000; a3 = 32'h00100000;  s = 10;
		#5 a0 = 32'hF1000000; a1 = 32'h01000000; a2 = 32'hF1000000; a3 = 32'h01000000;  s = 10;
		#5 a0 = 32'hF0000000; a1 = 32'h10000000; a2 = 32'hF0000000; a3 = 32'h10000000;  s = 10;
		#5 a0 = 32'hF00000BA; a1 = 32'h000000BA; a2 = 32'hF00000BA; a3 = 32'h000000BA;  s = 11;
		#5 a0 = 32'hF0000C00; a1 = 32'h00000C00; a2 = 32'hF0000C00; a3 = 32'h00000C00;  s = 11;
		#5 a0 = 32'hF000D000; a1 = 32'h0000D000; a2 = 32'hF000D000; a3 = 32'h0000D000;  s = 11;
		#5 a0 = 32'h00000000; a1 = 32'h00000000; a2 = 32'h00000000; a3 = 32'h00000000;  s = 11;
		#5 a0 = 32'h00000001; a1 = 32'h00000001; a2 = 32'h00000001; a3 = 32'h00000001;  s = 00;
		#5 a0 = 32'h00000010; a1 = 32'h00000010; a2 = 32'h00000010; a3 = 32'h00000010;  s = 00;
		#5 a0 = 32'h00000100; a1 = 32'h00000100; a2 = 32'h00000100; a3 = 32'h00000100;  s = 00;
		#5 a0 = 32'h00001000; a1 = 32'h00001000; a2 = 32'h00001000; a3 = 32'h00001000;  s = 00;
		#5 a0 = 32'h00010000; a1 = 32'h00010000; a2 = 32'h00010000; a3 = 32'h00010000;  s = 00;
		#5 a0 = 32'h00100000; a1 = 32'h00100000; a2 = 32'h00100000; a3 = 32'h00100000;  s = 00;
		#5 a0 = 32'h01000000; a1 = 32'h01000000; a2 = 32'h01000000; a3 = 32'h01000000;  s = 10;
		#5 a0 = 32'h10000000; a1 = 32'h10000000; a2 = 32'h10000000; a3 = 32'h10000000;  s = 10;
		#5 a0 = 32'h000000BA; a1 = 32'h000000BA; a2 = 32'h000000BA; a3 = 32'h000000BA;  s = 11;
		#5 a0 = 32'h00000C00; a1 = 32'h00000C00; a2 = 32'h00000C00; a3 = 32'h00000C00;  s = 11;
		#5 a0 = 32'h0000D000; a1 = 32'h0000D000; a2 = 32'h0000D000; a3 = 32'h0000D000;  s = 11;
	
	end
	
endmodule
