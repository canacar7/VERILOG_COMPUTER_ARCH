`timescale 1ns / 1ps
module islemler(a,b,x,y,z);
    input  [15:00] a;                                  // 16 bits
    input  [15:00] b;                                  // 16 bits
    output [31:07] x;                                  // sum high
    output [31:07] y;                                  // carry high
    output [06:00] z;                                  // sum low
    reg    [15:00] p [15:00];                          // p[i][j]
    parameter zero = 1'b0;                             // constant 0
    integer i, j;
    always @ * begin
        for (i = 0; i < 16; i = i + 1)
            for (j = 0; j < 16; j = j + 1)
                p[i][j] = a[i] & b[j];                 // p[i][j]=a[i]&b[j]
    end
    
     // level 1 ------------------------------------------------------------
    wire  [4:0] s1 [28:1]; //en fazla kullanÄ±an csa sayÄ±sÄ± 5 tane  
    wire  [4:0] c1 [29:2]; //level 1 icin sum ve carry tanimlari
    //     31:
    //     30:   p[15][15]
    //     29:   p[14][15] , p[15][14]
    csa a1_28_0 (p[13][15] , p[14][14] , p[15][13], s1[28][0], c1[29][0]);
    csa a1_27_0 (p[12][15] , p[13][14] , p[14][13], s1[27][0], c1[28][0]);
    //     27:   p[15][12] 
    csa a1_26_1 (p[11][15] , p[12][14] , p[13][13], s1[26][1], c1[27][1]);
    csa a1_26_0 (p[14][12] , p[15][11] , zero     , s1[26][0], c1[27][0]);
    csa a1_25_1 (p[10][15] , p[11][14] , p[12][13], s1[25][1], c1[26][1]);
    csa a1_25_0 (p[13][12] , p[14][11] , p[15][10], s1[25][0], c1[26][0]);
    csa a1_24_1 (p[9][15]  , p[10][14] , p[11][13], s1[24][1], c1[25][1]);
    csa a1_24_0 (p[12][12] , p[13][11] , p[14][10], s1[24][0], c1[25][0]);
    //     24:   p[15][9] 
    csa a1_23_2 (p[8][15]  ,p[9][14]   , p[10][13] , s1[23][2], c1[24][2]);
    csa a1_23_1 (p[11][12] ,p[12][11]  , p[13][10] , s1[23][1], c1[24][1]);
    csa a1_23_0 (p[14][9]  ,p[15][8]   , zero      , s1[23][0], c1[24][0]);
    csa a1_22_2 (p[7][15]  ,p[8][14]   , p[9][13]  , s1[22][2], c1[23][2]);
    csa a1_22_1 (p[10][12] ,p[11][11]  , p[12][10] , s1[22][1], c1[23][1]);
    csa a1_22_0 (p[13][9]  ,p[14][8]   , p[15][7]  , s1[22][0], c1[23][0]);
    csa a1_21_2 (p[6][15]  ,p[7][14]   , p[8][13]  , s1[21][2], c1[22][2]);
    csa a1_21_1 (p[9][10]  ,p[10][11]  , p[11][10] , s1[21][1], c1[22][1]);
    csa a1_21_0 (p[12][9]  ,p[13][8]   , p[14][7]  , s1[21][0], c1[22][0]);
    //     21:   p[15][6]
    csa a1_20_3 (p[5][15]  ,p[6][14]   , p[7][13]  , s1[20][3], c1[21][3]);
    csa a1_20_2 (p[8][12]  ,p[9][11]   , p[10][10] , s1[20][2], c1[21][2]);
    csa a1_20_1 (p[11][9]  ,p[12][8]   , p[13][7]  , s1[20][1], c1[21][1]);
    csa a1_20_0 (p[14][6]  ,p[15][5]   , zero      , s1[20][0], c1[21][0]);
    csa a1_19_3 (p[4][15]  ,p[5][14]   , p[6][13]  , s1[19][3], c1[20][3]);
    csa a1_19_2 (p[7][12]  ,p[8][11]   , p[9][10]  , s1[19][2], c1[20][2]);
    csa a1_19_1 (p[10][9]  ,p[11][8]   , p[12][7]  , s1[19][1], c1[20][1]);
    csa a1_19_0 (p[13][6]  ,p[14][5]   , p[15][4]  , s1[19][0], c1[20][0]); 
    csa a1_18_3 (p[3][15]  ,p[4][14]   , p[5][13]  , s1[18][3], c1[19][3]);
    csa a1_18_2 (p[6][12]  ,p[7][11]   , p[8][10]  , s1[18][2], c1[19][2]);
    csa a1_18_1 (p[9][9]  ,p[10][8]    , p[11][7]  , s1[18][1], c1[19][1]);
    csa a1_18_0 (p[12][6]  ,p[13][5]   , p[14][4]  , s1[18][0], c1[19][0]); 
    //     18:   p[15][3]
    csa a1_17_4 (p[2][15]  ,p[3][14]   , p[4][13]  , s1[17][4], c1[18][4]);
    csa a1_17_3 (p[5][12]  ,p[6][11]   , p[7][10]  , s1[17][3], c1[18][3]);
    csa a1_17_2 (p[8][9]   ,p[9][8]    , p[10][7]  , s1[17][2], c1[18][2]);
    csa a1_17_1 (p[11][6]  ,p[12][5]   , p[13][4]  , s1[17][1], c1[18][1]);
    csa a1_17_0 (p[14][3]  ,p[15][2]   , zero      , s1[17][0], c1[18][0]);
    csa a1_16_4 (p[1][15]  ,p[2][14]   , p[3][13]  , s1[16][4], c1[17][4]);
    csa a1_16_3 (p[4][12]  ,p[5][11]   , p[6][10]  , s1[16][3], c1[17][3]);
    csa a1_16_2 (p[7][9]   ,p[8][8]    , p[9][7]   , s1[16][2], c1[17][2]);
    csa a1_16_1 (p[10][6]  ,p[11][5]   , p[12][4]  , s1[16][1], c1[17][1]);
    csa a1_16_0 (p[13][3]  ,p[14][2]   , p[15][1]  , s1[16][0], c1[17][0]);
    csa a1_15_4 (p[0][15]  ,p[1][14]   , p[2][13]  , s1[15][4], c1[16][4]);
    csa a1_15_3 (p[3][12]  ,p[4][11]   , p[5][10]  , s1[15][3], c1[16][3]);
    csa a1_15_2 (p[6][9]   ,p[7][8]    , p[8][7]   , s1[15][2], c1[16][2]);
    csa a1_15_1 (p[9][6]   ,p[10][5]   , p[11][4]  , s1[15][1], c1[16][1]);
    csa a1_15_0 (p[12][3]  ,p[13][2]   , p[14][1]  , s1[15][0], c1[16][0]);
    //     15:   p[15][0]
    csa a1_14_4 (p[0][14]  ,p[1][13]   , p[2][12]  , s1[14][4], c1[15][4]);
    csa a1_14_3 (p[3][11]  ,p[4][10]   , p[5][9]   , s1[14][3], c1[15][3]);
    csa a1_14_2 (p[6][8]   ,p[7][7]    , p[8][6]   , s1[14][2], c1[15][2]);
    csa a1_14_1 (p[9][5]   ,p[10][4]   , p[11][3]  , s1[14][1], c1[15][1]);
    csa a1_14_0 (p[12][2]  ,p[13][1]   , p[14][0]  , s1[14][0], c1[15][0]);
    csa a1_13_4 (p[0][13]  ,p[1][12]   , p[2][11]  , s1[13][4], c1[14][4]);
    csa a1_13_3 (p[3][10]  ,p[4][9]    , p[5][8]   , s1[13][3], c1[14][3]);
    csa a1_13_2 (p[6][7]   ,p[7][6]    , p[8][5]   , s1[13][2], c1[14][2]);
    csa a1_13_1 (p[9][4]   ,p[10][3]   , p[11][2]  , s1[13][1], c1[14][1]);
    csa a1_13_0 (p[12][1]  ,p[13][0]   , zero      , s1[13][0], c1[14][0]);
    csa a1_12_3 (p[0][12]  ,p[1][11]   , p[2][10]  , s1[12][3], c1[13][3]);
    csa a1_12_2 (p[3][9]   ,p[4][8]    , p[5][7]   , s1[12][2], c1[13][2]);
    csa a1_12_1 (p[6][6]   ,p[7][5]    , p[8][4]   , s1[12][1], c1[13][1]);
    csa a1_12_0 (p[9][3]   ,p[10][2]   , p[11][1]  , s1[12][0], c1[13][0]);
    //     12:   p[12][0] 
    csa a1_11_3 (p[0][11]  ,p[1][10]   , p[2][9]   , s1[11][3], c1[12][3]);
    csa a1_11_2 (p[3][8]   ,p[4][7]    , p[5][6]   , s1[11][2], c1[12][2]);
    csa a1_11_1 (p[6][5]   ,p[7][4]    , p[8][3]   , s1[11][1], c1[12][1]);
    csa a1_11_0 (p[9][2]   ,p[10][1]   , p[11][0]  , s1[11][0], c1[12][0]);
    csa a1_10_3 (p[0][10]  ,p[1][9]    , p[2][8]   , s1[10][3], c1[11][3]);
    csa a1_10_2 (p[3][7]   ,p[4][6]    , p[5][5]   , s1[10][2], c1[11][2]);
    csa a1_10_1 (p[6][4]   ,p[7][3]    , p[8][2]   , s1[10][1], c1[11][1]);
    csa a1_10_0 (p[9][1]   ,p[10][0]   , zero      , s1[10][0], c1[11][0]);
    csa a1_9_2  (p[0][9]   ,p[1][8]    , p[2][7]   , s1[9][2] ,  c1[10][2]);
    csa a1_9_1  (p[3][6]   ,p[4][5]    , p[5][4]   , s1[9][1] ,  c1[10][1]);
    csa a1_9_0  (p[6][3]   ,p[7][2]    , p[8][1]   , s1[9][0] ,  c1[10][0]);
   //      9:    p[9][0] 
    csa a1_8_2  (p[0][8]   ,p[1][7]    , p[2][6]   , s1[8][2] ,  c1[9][2]);
    csa a1_8_1  (p[3][5]   ,p[4][4]    , p[5][3]   , s1[8][1] ,  c1[9][1]);
    csa a1_8_0  (p[6][2]   ,p[7][1]    , p[8][0]   , s1[8][0] ,  c1[9][0]);  
    csa a1_7_2  (p[0][7]   ,p[1][6]    , p[2][5]   , s1[7][2] ,  c1[8][2]);
    csa a1_7_1  (p[3][4]   ,p[4][3]    , p[5][2]   , s1[7][1] ,  c1[8][1]);
    csa a1_7_0  (p[6][1]   ,p[7][0]    , zero      , s1[7][0] ,  c1[8][0]); 
    csa a1_6_1  (p[0][6]   ,p[1][5]    , p[2][4]   , s1[6][1] ,  c1[7][1]);
    csa a1_6_0  (p[3][3]   ,p[4][2]    , p[5][1]   , s1[6][0] ,  c1[7][0]); 
    //      6:   p[6][0]
    csa a1_5_1  (p[0][5]   ,p[1][4]    , p[2][3]   , s1[5][1] ,  c1[6][1]);
    csa a1_5_0  (p[3][2]   ,p[4][1]    , p[5][0]   , s1[5][0] ,  c1[6][0]);
    csa a1_4_1  (p[0][4]   ,p[1][3]    , p[2][2]   , s1[4][1] ,  c1[5][1]);
    csa a1_4_0  (p[3][1]   ,p[4][0]    , zero      , s1[4][0] ,  c1[5][0]);
    csa a1_3_0  (p[0][3]   ,p[1][2]    , p[2][1]   , s1[3][0] ,  c1[4][0]); 
    //      3:   p[3][0]
    csa a1_2_0  (p[0][2]   ,p[1][1]    , p[2][0]   , s1[2][0] ,  c1[3][0]); 
    csa a1_1_0  (p[0][1]   ,p[0][1]    , zero      , s1[1][0] ,  c1[2][0]); 
    //     0:   p[0][0]
// level 2 ------------------------------------------------------------    
    wire  [3:0] s2 [29:2];
    wire  [3:0] c2 [30:3];
    //     31:
    //     30:   p[15][15]
    csa a2_29_0 (p[14][15], p[15][14], c1[29][0], s2[29][0], c2[30][0]);
    csa a2_28_0 (s1[28][0], c1[28][0], zero     , s2[28][0], c2[29][0]);
    csa a2_27_0 (s1[27][0], p[15][12], c1[27][1], s2[27][0], c2[28][0]);
    //     27:   c1[27][0]
    csa a2_26_0 (s1[26][1], s1[26][0], c1[26][1], s2[26][0], c2[27][0]);
    //     26:   c1[26][0]
    csa a2_25_0 (s1[25][1], s1[25][0], c1[25][1], s2[25][0], c2[26][0]);
    //     25:   c1[25][0]
    csa a2_24_1 (s1[24][1], s1[24][0], p[15][9] , s2[24][1], c2[25][1]);
    csa a2_24_0 (c1[24][2], c1[24][1], c1[24][0], s2[24][0], c2[25][0]);
    csa a2_23_1 (s1[23][2], s1[23][1], s1[23][0], s2[23][1], c2[24][1]);
    csa a2_23_0 (c1[23][2], c1[23][1], c1[23][0], s2[23][0], c2[24][0]);
    csa a2_22_1 (s1[22][2], s1[22][1], s1[22][0], s2[22][1], c2[23][1]);
    csa a2_22_0 (c1[22][2], c1[22][1], c1[22][0], s2[22][0], c2[23][0]);
    csa a2_21_2 (s1[21][2], s1[21][1], s1[21][0], s2[21][2], c2[22][2]);
    csa a2_21_1 (p[15][6] , c1[21][3], c1[21][2], s2[21][1], c2[22][1]);
    csa a2_21_0 (c1[21][1], c1[21][0],      zero, s2[21][0], c2[22][0]);
    csa a2_20_2 (s1[20][3], s1[20][2], s1[20][1], s2[20][2], c2[21][2]);
    csa a2_20_1 (s1[20][0], c1[20][3], c1[20][2], s2[20][1], c2[21][1]);
    csa a2_20_0 (c1[20][1], c1[20][0],      zero, s2[20][0], c2[21][0]);
    csa a2_19_2 (s1[19][3], s1[19][2], s1[19][1], s2[19][2], c2[20][2]);
    csa a2_19_1 (s1[19][0], c1[19][3], c1[19][2], s2[19][1], c2[20][1]);
    csa a2_19_0 (c1[19][1], c1[19][0],      zero, s2[19][0], c2[20][0]);
    csa a2_18_2 (s1[18][3], s1[18][2], s1[18][1], s2[18][2], c2[19][2]);
    csa a2_18_1 (s1[18][0], p[15][3] , c1[18][4], s2[18][1], c2[19][1]);
    csa a2_18_0 (c1[18][3], c1[18][2], c1[18][1], s2[18][0], c2[19][0]);
    //     18:   c1[18][0]
    csa a2_17_2 (s1[17][4], s1[17][3], s1[17][2], s2[17][2], c2[18][2]);
    csa a2_17_1 (s1[17][1], s1[17][0], c1[17][4], s2[17][1], c2[18][1]);
    csa a2_17_0 (c1[17][3], c1[17][2], c1[17][1], s2[17][0], c2[18][0]);
    //     17:   c1[17][0]
    csa a2_16_2 (s1[16][4], s1[16][3], s1[16][2], s2[16][2], c2[17][2]);
    csa a2_16_1 (s1[16][1], s1[16][0], c1[16][4], s2[16][1], c2[17][1]);
    csa a2_16_0 (c1[16][3], c1[16][2], c1[16][1], s2[16][0], c2[17][0]);
    //     16:   c1[16][0]
    csa a2_15_3 (s1[15][4], s1[15][3], s1[15][2] , s2[15][3], c2[16][3]);
    csa a2_15_2 (s1[15][1], s1[15][0], p[15][0]  , s2[15][2], c2[16][2]);
    csa a2_15_1 (c1[15][4], c1[15][3], c1[15][2] , s2[15][1], c2[16][1]);
    csa a2_15_0 (c1[15][1], c1[15][0],  zero     , s2[15][0], c2[16][0]);
    csa a2_14_2 (s1[14][4], s1[14][3], s1[14][2] , s2[14][2], c2[15][2]);
    csa a2_14_1 (s1[14][1], s1[14][0], c1[14][4] , s2[14][1], c2[15][1]);
    csa a2_14_0 (c1[14][3], c1[14][2], c1[14][1] , s2[14][0], c2[15][0]);
    //     14:   c1[14][0]
    csa a2_13_2 (s1[13][4], s1[13][3], s1[13][2] , s2[13][2], c2[14][2]);
    csa a2_13_1 (s1[13][1], s1[13][0], c1[13][3] , s2[13][1], c2[14][1]);
    csa a2_13_0 (c1[13][2], c1[13][1], c1[13][0] , s2[13][0], c2[14][0]);
    csa a2_12_2 (s1[12][3], s1[12][2], s1[12][1] , s2[12][2], c2[13][2]);
    csa a2_12_1 (s1[12][0], p[12][0] , c1[12][3] , s2[12][1], c2[13][1]);
    csa a2_12_0 (c1[12][2], c1[12][1], c1[12][0] , s2[12][0], c2[13][0]);
    csa a2_11_2 (s1[11][3], s1[11][2], s1[11][1] , s2[11][2], c2[12][2]);
    csa a2_11_1 (s1[11][0], c1[11][3], c1[11][2] , s2[11][1], c2[12][1]);
    csa a2_11_0 (c1[11][1], c1[11][0], zero      , s2[11][0], c2[12][0]);
    csa a2_10_1 (s1[10][3], s1[10][2], s1[10][1] , s2[10][1], c2[11][1]);
    csa a2_10_0 (s1[10][0], c1[10][2], c1[10][1] , s2[10][0], c2[11][0]);
    //     10:   c1[10][0]
    csa a2_9_1  (s1[9][2] , s1[9][1], s1[9][0]   , s2[9][1], c2[10][1]);
    csa a2_9_0  (p[9][0]  , c1[9][2], c1[9][1]   , s2[9][0], c2[10][0]);
    //     9:   c1[9][0]
    csa a2_8_1  (s1[8][2] , s1[8][1], s1[8][0]   , s2[8][1], c2[9][1]);
    csa a2_8_0  (c1[8][1] , c1[8][0], c1[8][0]   , s2[8][0], c2[9][0]);
    csa a2_7_1  (s1[7][2] , s1[7][1], s1[7][0]   , s2[7][1], c2[8][1]);
    csa a2_7_0  (c1[7][1] , c1[7][0], zero       , s2[7][0], c2[8][0]);
    csa a2_6_1 (s1[6][1]  , s1[6][0], p[6][0]    , s2[6][1], c2[7][1]);
    csa a2_6_0 (c1[6][1]  , c1[6][0],      zero  , s2[6][0], c2[7][0]);
    csa a2_5_0 (s1[5][1]  , s1[5][0], c1[5][1]  , s2[5][0], c2[6][0]);
    //     5:   c1[5][0]
    csa a2_4_0 (s1[4][1], s1[4][0], c1[4][0]  , s2[4][0], c2[5][0]);
    csa a2_3_0 (s1[3][0], p[3][0]  , c1[3][0]  , s2[3][0], c2[4][0]);
    csa a2_2_0 (s1[2][0], c1[2][0],     zero  , s2[2][0], c2[3][0]);
    //    1:   s1[1][0]
    //    0:   p[0][0]
    
// level 3 ------------------------------------------------------------     
    wire  [2:0] s3 [30:3];
    wire  [2:0] c3 [31:4];
    //     31:
    csa a3_30_0 (p[15][15] , c2[30][0],       zero, s3[30][0], c3[31][0]);
    csa a3_29_0 (s2[29][0] , c2[29][0],       zero, s3[29][0], c3[30][0]);
    csa a3_28_0 (s2[28][0] , c2[28][0],       zero, s3[28][0], c3[29][0]);
    csa a3_27_0 (s2[27][0] , c1[27][0],  c2[27][0], s3[27][0], c3[28][0]);
    csa a3_26_0 (s2[26][0] , c1[26][0],  c2[26][0], s3[26][0], c3[27][0]);
    csa a3_25_0 (s2[25][0] , c1[25][0],  c2[25][1], s3[25][0], c3[26][0]);
    //     25:   c2[25][0]
    csa a3_24_0 (s2[24][1] , s2[24][0],  c2[24][1], s3[24][0], c3[25][0]);
    //     24:   c2[24][0]
    csa a3_23_0 (s2[23][1] , s2[23][0],  c2[23][1], s3[23][0], c3[24][0]);
    //     23:   c2[23][0]
    csa a3_22_1 (s2[22][1] , s2[22][0],  c2[22][2]     , s3[22][1], c3[23][1]);
    csa a3_22_0 (c2[22][1] , c2[22][0],  zero          , s3[22][0], c3[23][0]);
    csa a3_21_1 (s2[21][2] , s2[21][1],  s2[21][0]     , s3[21][1], c3[22][1]);
    csa a3_21_0 (c2[21][2] , c2[21][1],  c2[21][0]     , s3[21][0], c3[22][0]);
    csa a3_20_1 (s2[20][2] , s2[20][1],  s2[20][0]     , s3[20][1], c3[21][1]);
    csa a3_20_0 (c2[20][2] , c2[20][1],  c2[20][0]     , s3[20][0], c3[21][0]);
    csa a3_19_1 (s2[19][2] , s2[19][1],  s2[19][0]     , s3[19][1], c3[20][1]);
    csa a3_19_0 (c2[19][2] , c2[19][1],  c2[19][0]     , s3[19][0], c3[20][0]);    
    csa a3_18_1 (s2[18][2] , s2[18][1],  s2[18][0]     , s3[18][1], c3[19][1]);
    csa a3_18_0 (c1[18][0] ,c2[18][2] ,  c2[18][1]     , s3[18][0], c3[19][0]); 
    //          c2[18][0]
    csa a3_17_1 (s2[17][2] , s2[17][1],  s2[17][0]     , s3[17][1], c3[18][1]);
    csa a3_17_0 (c1[17][0] , c2[17][2] ,  c2[17][1]    , s3[17][0], c3[18][0]); 
    //          c2[17][0]  
    csa a3_16_2 (s2[16][2] , s2[16][1],  s2[16][0]     , s3[16][2], c3[17][2]);
    csa a3_16_1 (c1[16][0] , c2[16][3],  c2[16][2]     , s3[16][1], c3[17][1]); 
    csa a3_16_0 (c2[16][1] , c2[16][0],  zero          , s3[16][0], c3[17][0]); 
    csa a3_15_1 (s2[15][3] , s2[15][2],  s2[15][1]     , s3[15][1], c3[16][1]);
    csa a3_15_0 (s2[15][0] , c2[15][2],  c2[15][1]     , s3[15][0], c3[16][0]);
    //          c2[15][0]
    csa a3_14_1 (s2[14][2] , s2[14][1],  s2[14][0]     , s3[14][1], c3[15][1]);
    csa a3_14_0 (c1[14][0] , c2[14][2],  s2[14][1]     , s3[14][0], c3[15][0]);
    //          c2[14][0]    
    csa a3_13_1 (s2[13][2] , s2[13][1],  s2[13][0]     , s3[13][1], c3[14][1]);
    csa a3_13_0 (c2[13][2] , c2[13][1],  c2[13][0]     , s3[13][0], c3[14][0]);
    csa a3_12_1 (s2[12][2] , s2[12][1],  s2[12][0]     , s3[12][1], c3[13][1]);
    csa a3_12_0 (c2[12][2] , c2[12][1],  c2[12][0]     , s3[12][0], c3[13][0]);
    csa a3_11_1 (s2[11][2] , s2[11][1],  s2[11][0]     , s3[11][1], c3[12][1]);
    csa a3_11_0 (c2[11][1] , c2[11][0],  zero          , s3[11][0], c3[12][0]);
    csa a3_10_1 (s2[10][1] , s2[10][0],  c1[10][0]     , s3[10][1], c3[11][1]);
    csa a3_10_0 (c2[10][1] , c2[10][0],  zero          , s3[10][0], c3[11][0]);
    csa a3_09_1 (s2[9][1], s2[9][0]   ,  c1[9][0]      , s3[9][1], c3[10][1]);
    csa a3_09_0 (c2[9][1], c2[9][0]   ,      zero      , s3[9][0], c3[10][0]);
    csa a3_08_0 (s2[8][1], s2[8][0]   , c2[8][1]      , s3[8][0], c3[9][0]);
    //     08:   c2[8][0]
    csa a3_07_0 (s2[7][1], s2[7][0]   , c2[7][1]      , s3[7][0], c3[8][0]);
    //     07:   c[7][0]
    csa a3_06_0 (s2[6][1], s2[6][0]   , c2[6][0]      , s3[6][0], c3[7][0]);
    csa a3_05_0 (s2[5][0], c1[5][0]   , c2[5][0]      , s3[5][0], c3[6][0]);
    csa a3_04_0 (s2[4][0], c2[4][0]   ,      zero      , s3[4][0], c3[5][0]);
    csa a3_03_0 (s2[3][0], c2[3][0]   ,      zero      , s3[3][0], c3[4][0]);
    //     02:   s2[2][0]
    //     01:   s1[1][0]
    //     00:   p[0][0]
    
     // level 4 ------------------------------------------------------------
    wire  [1:0] s4 [30:4];
    wire  [1:0] c4 [31:5];
    
       
     //     31:   c3[31][0]
    csa a4_30_0 (s3[30][0], c3[30][0],      zero, s4[30][0], c4[31][0]);
    csa a4_29_0 (s3[29][0], c3[29][0],      zero, s4[29][0], c4[30][0]);
    csa a4_28_0 (s3[28][0], c3[28][0],      zero, s4[28][0], c4[29][0]);
    csa a4_27_0 (s3[27][0], c3[27][0],      zero, s4[27][0], c4[28][0]);
    csa a4_26_0 (s3[26][0], c3[26][0],      zero, s4[26][0], c4[27][0]);
    csa a4_25_0 (s3[25][0], c2[25][0], c3[25][0], s4[25][0], c4[26][0]);
    csa a4_24_0 (s3[24][0], c2[24][0], c3[24][0], s4[24][0], c4[25][0]);
    csa a4_23_0 (s3[23][0], c2[23][0], c3[23][1], s4[23][0], c4[24][0]);
    //     23:   c3[23][0]
    csa a4_22_0 (s3[22][1], s3[22][0], c3[22][1], s4[22][0], c4[23][0]);
    //     22:   c3[22][0          
    csa a4_21_0 (s3[21][1], s3[21][0], c3[21][1], s4[21][0], c4[22][0]);
    //     21:   c3[21][0]         
    csa a4_20_0 (s3[20][1], s3[20][0], c3[20][1], s4[20][0], c4[21][0]);
    //     20:   c3[20][0]         
    csa a4_19_0 (s3[19][1], s3[19][0], c3[19][1], s4[19][0], c4[20][0]);
    //     19:   c3[19][0]         
    csa a4_18_1 (s3[18][1], s3[18][0], c2[18][0], s4[18][1], c4[19][1]);
    csa a4_18_0 (c3[18][1], c3[18][0], zero     , s4[18][0], c4[19][0]);
    csa a4_17_1 (s3[17][1], s3[17][0], c2[17][0], s4[17][1], c4[18][1]);
    csa a4_17_0 (c3[17][2], c3[17][1], c3[17][0], s4[17][0], c4[18][0]);     
    csa a4_16_1 (s3[16][2], s3[16][1], s3[16][0], s4[16][1], c4[17][1]);
    csa a4_16_0 (c3[16][1], c3[16][0], zero     , s4[16][0], c4[17][0]); 
    csa a4_15_1 (s3[15][1], s3[15][0], c2[15][0], s4[15][1], c4[16][1]);
    csa a4_15_0 (c3[15][1], c3[15][0], zero     , s4[15][0], c4[16][0]);
    csa a4_14_1 (s3[14][1], s3[14][0], c2[14][0], s4[14][1], c4[15][1]);
    csa a4_14_0 (c3[14][1], c3[14][0], zero     , s4[14][0], c4[15][0]);    
    csa a4_13_0 (s3[13][1], s3[13][0], c3[13][1], s4[13][0], c4[14][0]);
    //     13:   c3[13][0]    
    csa a4_12_0 (s3[12][1], s3[12][0], c3[12][1], s4[12][0], c4[13][0]);
    //     12:   c3[12][0]
    csa a4_11_0 (s3[11][1], s3[11][0], c3[11][1], s4[11][0], c4[12][0]);
    //     11:   c3[11][0]    
    csa a4_10_0 (s3[10][1], s3[10][0], c3[10][1], s4[10][0], c4[11][0]);
    //     10:   c3[10][0]
    csa a4_9_0 (s3[9][1], s3[9][0], c3[10][0],    s4[9][0], c4[10][0]);
    csa a4_8_0 (s3[8][0], c2[8][0], c3[8][0],     s4[8][0], c4[9][0]);
    csa a4_7_0 (s3[7][0], c2[7][0], c3[7][0],     s4[7][0], c4[8][0]);
    csa a4_6_0 (s3[6][0], c3[6][0], zero    ,     s4[6][0], c4[7][0]);
    csa a4_5_0 (s3[5][0], c3[5][0], zero    ,     s4[5][0], c4[6][0]);
    csa a4_4_0 (s3[4][0], c3[4][0], zero    ,     s4[4][0], c4[5][0]);
    //     03:   s3[3][0]
    //     02:   s2[2][0]
    //     01:   s1[1][0]
    //     00:   p[0][0]
   
   
   // level 5 ------------------------------------------------------------
    wire  [0:0] s5 [31:5];
    wire  [0:0] c5 [32:6];
    
    
    csa a5_31_0 (c3[31][0], c4[31][0],      zero, s5[31][0], c5[32][0]);
    csa a5_30_0 (s4[30][0], c4[30][0],      zero, s5[30][0], c5[31][0]);
    csa a5_29_0 (s4[29][0], c4[29][0],      zero, s5[29][0], c5[30][0]);
    csa a5_28_0 (s4[28][0], c4[28][0],      zero, s5[28][0], c5[29][0]);
    csa a5_27_0 (s4[27][0], c4[27][0],      zero, s5[27][0], c5[28][0]);
    csa a5_26_0 (s4[26][0], c4[26][0],      zero, s5[26][0], c5[27][0]);
    csa a5_25_0 (s4[25][0], c4[25][0],      zero, s5[25][0], c5[26][0]);
    csa a5_24_0 (s4[24][0], c4[24][0],      zero, s5[24][0], c5[25][0]);
    csa a5_23_0 (s4[23][0], c3[23][0], c4[23][0], s5[23][0], c5[24][0]);
    csa a5_22_0 (s4[22][0], c3[22][0], c4[22][0], s5[22][0], c5[23][0]);
    csa a5_21_0 (s4[21][0], c3[21][0], c4[21][0], s5[21][0], c5[22][0]);
    csa a5_20_0 (s4[20][0], c3[20][0], c4[20][0], s5[20][0], c5[21][0]);
    csa a5_19_0 (s4[19][0], c3[19][0], c4[19][1], s5[19][0], c5[20][0]);
    //     19:   c4[19][0]
    csa a5_18_0 (s4[18][1], s4[18][0], c4[18][1], s5[18][0], c5[19][0]);
    //     18:   c4[18][0]
    csa a5_17_0 (s4[17][1], s4[17][0], c4[17][1], s5[17][0], c5[18][0]);
    //     17:   c4[17][0] 
    csa a5_16_0 (s4[16][1], s4[16][0], c4[16][1], s5[16][0], c5[17][0]);
    //     16:   c4[16][0] 
    csa a5_15_0 (s4[15][1], s4[15][0], c4[15][1], s5[15][0], c5[16][0]);
    //     15:   c4[15][0]
    csa a5_14_0 (s4[14][1], s4[14][0], c4[14][0], s5[14][0], c5[15][0]);
    csa a5_13_0 (s4[13][0], c3[13][0], c4[13][0], s5[13][0], c5[14][0]);
    csa a5_12_0 (s4[12][0], c3[12][0], c4[12][0], s5[12][0], c5[13][0]);
    csa a5_11_0 (s4[11][0], c3[11][0], c4[11][0], s5[11][0], c5[12][0]);
    csa a5_10_0 (s4[10][0], c3[10][0], c4[10][0], s5[10][0], c5[11][0]);
    csa a5_9_0  (s4[9][0] , c4[9][0] , zero     , s5[9][0] , c5[10][0]);
    csa a5_8_0  (s4[8][0] , c4[8][0] , zero     , s5[8][0] , c5[9][0]);
    csa a5_7_0  (s4[7][0] , c4[7][0] , zero     , s5[7][0] , c5[8][0]);
    csa a5_6_0  (s4[6][0] , c4[6][0] , zero     , s5[6][0] , c5[7][0]);
    csa a5_5_0  (s4[5][0] , c4[5][0] , zero     , s5[5][0] , c5[6][0]);
    //     4:   s4[4][0]
    //     3:   s3[3][0]
    //     2:   s2[2][0]
    //     1:   s1[1][0]
    //     0:   p[0][0]

    // level 6 ------------------------------------------------------------
    wire  [0:0] s6 [31:6];
    wire  [0:0] c6 [32:7];
    
    csa a6_31_0 (s5[31][0], c5[31][0],      zero, s6[31][0], c6[32][0]);
    csa a6_30_0 (s5[30][0], c5[30][0],      zero, s6[30][0], c6[31][0]);
    csa a6_29_0 (s5[29][0], c5[29][0],      zero, s6[29][0], c6[30][0]);
    csa a6_28_0 (s5[28][0], c5[28][0],      zero, s6[28][0], c6[29][0]);
    csa a6_27_0 (s5[27][0], c5[27][0],      zero, s6[27][0], c6[28][0]);
    csa a6_26_0 (s5[26][0], c5[26][0],      zero, s6[26][0], c6[27][0]);
    csa a6_25_0 (s5[25][0], c5[25][0],      zero, s6[25][0], c6[26][0]);
    csa a6_24_0 (s5[24][0], c5[24][0],      zero, s6[24][0], c6[25][0]);
    csa a6_23_0 (s5[23][0], c5[23][0],      zero, s6[23][0], c6[24][0]);
    csa a6_22_0 (s5[22][0], c5[22][0],      zero, s6[22][0], c6[23][0]);
    csa a6_21_0 (s5[21][0], c5[21][0],      zero, s6[21][0], c6[22][0]);
    csa a6_20_0 (s5[20][0], c5[20][0],      zero, s6[20][0], c6[21][0]);
    csa a6_19_0 (s5[19][0], c4[19][0], c5[19][0], s6[19][0], c6[20][0]);
    csa a6_18_0 (s5[18][0], c4[18][0], c5[18][0], s6[18][0], c6[19][0]);
    csa a6_17_0 (s5[17][0], c4[17][0], c5[17][0], s6[17][0], c6[18][0]);
    csa a6_16_0 (s5[16][0], c4[16][0], c5[16][0], s6[16][0], c6[17][0]);
    csa a6_15_0 (s5[15][0], c4[15][0], c5[15][0], s6[15][0], c6[16][0]);
    csa a6_14_0 (s5[14][0], c5[14][0],      zero, s6[14][0], c6[15][0]);
    csa a6_13_0 (s5[13][0], c5[13][0],      zero, s6[13][0], c6[14][0]);
    csa a6_12_0 (s5[12][0], c5[12][0],      zero, s6[12][0], c6[13][0]);
    csa a6_11_0 (s5[11][0], c5[11][0],      zero, s6[11][0], c6[12][0]);
    csa a6_10_0 (s5[10][0], c5[10][0],      zero, s6[10][0], c6[11][0]);
    csa a6_9_0 (s5[09][0] , c5[09][0],      zero, s6[09][0], c6[10][0]);
    csa a6_8_0 (s5[08][0] , c5[08][0],      zero, s6[08][0], c6[09][0]);
    csa a6_7_0 (s5[07][0] , c5[07][0],      zero, s6[07][0], c6[08][0]);
    csa a6_6_0 (s5[06][0] , c5[06][0],      zero, s6[06][0], c6[07][0]);
    //     5:   s5[5][0]
    //     4:   s4[4][0]
    //     3:   s3[3][0]
    //     2:   s2[2][0]
    //     1:   s1[1][0]
    //     0:   p[0][0]
    
    
    assign x[31] = s6[31][0];                  assign y[31] = c6[31][0];
    assign x[30] = s6[30][0];                  assign y[30] = c6[30][0];
    assign x[29] = s6[29][0];                  assign y[29] = c6[29][0];
    assign x[28] = s6[28][0];                  assign y[28] = c6[28][0];
    assign x[27] = s6[27][0];                  assign y[27] = c6[27][0];
    assign x[26] = s6[26][0];                  assign y[26] = c6[26][0];
    assign x[25] = s6[25][0];                  assign y[25] = c6[25][0];
    assign x[24] = s6[24][0];                  assign y[24] = c6[24][0];
    assign x[23] = s6[23][0];                  assign y[23] = c6[23][0];
    assign x[22] = s6[22][0];                  assign y[22] = c6[22][0];
    assign x[21] = s6[21][0];                  assign y[21] = c6[21][0];
    assign x[20] = s6[20][0];                  assign y[20] = c6[20][0];
    assign x[19] = s6[19][0];                  assign y[19] = c6[19][0];
    assign x[18] = s6[18][0];                  assign y[18] = c6[18][0];
    assign x[17] = s6[17][0];                  assign y[17] = c6[17][0];
    assign x[16] = s6[16][0];                  assign y[16] = c6[16][0];
    assign x[15] = s6[15][0];                  assign y[15] = c6[15][0];
    assign x[14] = s6[14][0];                  assign y[14] = c6[14][0];
    assign x[13] = s6[13][0];                  assign y[13] = c6[13][0];
    assign x[12] = s6[12][0];                  assign y[12] = c6[12][0];
    assign x[11] = s6[11][0];                  assign y[11] = c6[11][0];
    assign x[10] = s6[10][0];                  assign y[10] = c6[10][0];
    assign x[9]  = s6[9][0];                   assign y[9]  = c6[9][0];
    assign x[8]  = s6[8][0];                   assign y[8]  = c6[8][0];
    assign x[7]  = s6[7][0];                   assign y[7]  = c6[7][0];
    
    
    assign z[6] = s6[6][0];
    assign z[5] = s5[5][0];
    assign z[4] = s4[4][0];
    assign z[3] = s3[3][0];
    assign z[2] = s2[2][0];
    assign z[1] = s1[1][0];
    assign z[0] = p[0][0];
    
    
endmodule
