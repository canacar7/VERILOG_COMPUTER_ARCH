module odev64_bit(a,b,z,z_1,z_2,clk,rst);
    input   clk,rst;
    input   [31:0] a, b;                             // a, b
    output [63:0] z;                                // z = a * b
    output [63:0] z_1,z_2;
    reg     [31:0] abi[31:0];                         // a[i] & b[j]
    integer       i, j;
    reg  u;
	
	reg     [2 : 0] state, next_state;
	parameter       unsigned_durumu = 1'b0,
					signed_durumu   = 1'b1;
	

					
	always @(posedge clk or negedge rst) begin
		 if (rst) begin
			state <= signed_durumu;
		 end else 
			state <= next_state;
	end		

	always @(*) begin
		case(state)	
		
			unsigned_durumu : begin
                    for (j = 0; j < 32; j = j + 1)
                     for (i = 0; i < 32; i = i + 1)
                         abi[i][j] = a[i] & b[j];            
			    		next_state <= signed_durumu;
			    		u <= 1'b0;
				end
			 
							  
			signed_durumu : begin
					for (i = 0; i < 31; i = i + 1)
						for (j = 0; j < 31; j = j + 1)
							abi[i][j] = a[i] & b[j];           
					for (i = 0; i < 31; i = i + 1)
						abi[i][31] = ~(a[i] & b[31]);             
					for (j = 0; j < 31; j = j + 1)
						abi[31][j] = ~(a[31] & b[j]);             
					abi[31][31] = a[31] & b[31];
					next_state <= unsigned_durumu;
					u <= 1'b1;
	          end		
		endcase				  
    end
    
	assign z_1 = (({32'b0, abi[0][31:0]}              +        
                 {31'b0,   abi[1][31:0] ,  1'b0})      +        
                ({30'b0,   abi[2][31:0] ,  2'b0}       +        
                 {29'b0,   abi[3][31:0] ,  3'b0}))     +        
               (({28'b0,   abi[4][31:0] ,  4'b0}       +        
                 {27'b0,   abi[5][31:0] ,  5'b0})      +       
                ({26'b0,   abi[6][31:0] ,  6'b0}       +        
                 {25'b0,   abi[7][31:0] ,  7'b0}))     +         
               (({24'b0,   abi[8][31:0] ,  8'b0}       +        
                 {23'b0,   abi[9][31:0] ,  9'b0})      +       
                ({22'b0,   abi[10][31:0],  10'b0}      +        
                 {21'b0,   abi[11][31:0],  11'b0}))	  +
               (({20'b0,   abi[12][31:0],  12'b0}      +        
                 {19'b0,   abi[13][31:0],  13'b0})     +       
                ({18'b0,   abi[14][31:0],  14'b0}      +        
                 {17'b0,   abi[15][31:0],  15'b0}))	  +				 
               (({16'b0,   abi[16][31:0],  16'b0}      +        
                 {15'b0,   abi[17][31:0],  17'b0})     +       
                ({14'b0,   abi[18][31:0],  18'b0}      +        
                 {13'b0,   abi[19][31:0],  19'b0}))	  +	
               (({12'b0,   abi[20][31:0],  20'b0}      +        
                 {11'b0,   abi[21][31:0],  21'b0})     +       
                ({10'b0,   abi[22][31:0],  22'b0}      +        
                 {9'b0,    abi[23][31:0],  23'b0}))	  +				 
               (({8'b0,    abi[24][31:0],  24'b0}     +        
                 {7'b0,    abi[25][31:0],  25'b0})    +       
                ({6'b0,    abi[26][31:0],  26'b0}     +        
                 {5'b0,    abi[27][31:0],  27'b0}))   +				 
               (({4'b0,    abi[28][31:0],  28'b0}     +        
                 {3'b0,    abi[29][31:0],  29'b0})    +       
                ({2'b0,    abi[30][31:0],  30'b0}     +        
                 {1'b0,    abi[31][31:0],  31'b0}));				 
			 
	assign z_2 = (({32'b1, abi[0][31:0]}              +        
                 {31'b0,   abi[1][31:0] ,  1'b0})      +        
                ({30'b0,   abi[2][31:0] ,  2'b0}       +        
                 {29'b0,   abi[3][31:0] ,  3'b0}))     +        
               (({28'b0,   abi[4][31:0] ,  4'b0}       +        
                 {27'b0,   abi[5][31:0] ,  5'b0})      +       
                ({26'b0,   abi[6][31:0] ,  6'b0}       +        
                 {25'b0,   abi[7][31:0] ,  7'b0}))     +         
               (({24'b0,   abi[8][31:0] ,  8'b0}       +        
                 {23'b0,   abi[9][31:0] ,  9'b0})      +       
                ({22'b0,   abi[10][31:0],  10'b0}      +        
                 {21'b0,   abi[11][31:0],  11'b0}))	  +
               (({20'b0,   abi[12][31:0],  12'b0}      +        
                 {19'b0,   abi[13][31:0],  13'b0})     +       
                ({18'b0,   abi[14][31:0],  14'b0}      +        
                 {17'b0,   abi[15][31:0],  15'b0}))	  +				 
               (({16'b0,   abi[16][31:0],  16'b0}      +        
                 {15'b0,   abi[17][31:0],  17'b0})     +       
                ({14'b0,   abi[18][31:0],  18'b0}      +        
                 {13'b0,   abi[19][31:0],  19'b0}))	  +	
               (({12'b0,   abi[20][31:0],  20'b0}      +        
                 {11'b0,   abi[21][31:0],  21'b0})     +       
                ({10'b0,   abi[22][31:0],  22'b0}      +        
                 {9'b0,    abi[23][31:0],  23'b0}))	  +				 
               (({8'b0,    abi[24][31:0],  24'b0}     +        
                 {7'b0,    abi[25][31:0],  25'b0})    +       
                ({6'b0,    abi[26][31:0],  26'b0}     +        
                 {5'b0,    abi[27][31:0],  27'b0}))   +				 
               (({4'b0,    abi[28][31:0],  28'b0}     +        
                 {3'b0,    abi[29][31:0],  29'b0})    +       
                ({2'b0,    abi[30][31:0],  30'b0}     +        
                 {1'b1,    abi[31][31:0],  31'b0}));				 


     

    assign z = u ? z_2 : z_1;
endmodule
